`include "cpu.svh"

module cpu
    (
        input logic clk_100M, clk_en, rst,
        input logic [31:0] r_data,
        output logic wr_en,
        output logic [31:0] mem_addr, w_data,
        // debug addr/data and instr are for showing CPU information
        // on the FPGA (only useful in synthesis)
        input logic [4:0] rdbg_addr,
        output logic [31:0] rdbg_data,
        output logic [31:0] instr
    );
    // The CPU interfaces with main memory which is enabled by the
    // inputs and outputs of this module (r_data, wr_en, mem_addr, w_data)
    // You should create the register file, flip flops, and logic implementing
    // a simple datapath so that instructions can be loaded from main memory,
    // executed, and the results can be inspected in the register file, or in
    // main memory (once lw and sw are supported). You should also create a
    // control FSM that controls the behavior of the datapath depending on the
    // instruction that is currently executing. You may want to split the CPU
    // into one or more submodules.
    //
    // We have provided modules for you to use inside the CPU. Please see
    // the following files:
    // reg_file.sv (register file), reg_en.sv (register with enable and reset),
    // reg_reset.sv (register with only reset), alu.sv (ALU)
    // Useful constants and opcodes are provided in cpu.svh, which is included
    // at the top of this file.
    //
    // Place the instruction machine code (generated by your assembler, or the
    // provided assembler) in asm/instr.mem and it will be automatically
    // loaded into main memory starting at address 0x00400000. Make sure the memory
    // file is imported into Vivado first (`./tcl.sh refresh`).

    // PC logic
    logic [31:0] PC_prime, PC_real;

    // memory logic
    logic [31:0] Adr, RAM_out, Instr, Data;

    // instruction logic
    logic [5:0] opcode, funct;
    logic [4:0] rs, rt, rd, shamt;
    logic [15:0] imm;
    logic [25:0] addr;

    // register logic
    logic [4:0] Reg_A3;
    logic [31:0] Reg_WD3;
    logic [31:0] RD1_out, RD2_out, Reg_A, Reg_B;

    // ALU logic
    logic [31:0] SrcA, SrcB, SignImm, Zero, ALUResult, ALUOut, Shifted_2;

    // Jump logic
    logic [27:0] shifted_addr;
    logic [3:0] PC_first;
    logic [31:0] PCJump;

    // control signals
    logic IorD, MemWrite, IRWrite, PCWrite, Branch, ALUSrcA, RegWrite, PCEn, BNe;
    logic [3:0] ALUControl;
    logic [1:0] ALUSrcB, PCSrc, MemtoReg, RegDst;

    control control_unit (.*);
    assign wr_en = MemWrite;

        //PC update
        reg_en pc_update 
            (.clk(clk_100M), .en(PCEn), .d(PC_prime), .q(PC_real));
        // mux before RAM
        two_mux adress_mux 
            (.d_0(PC_real), .d_1(ALUOut), .z(Adr), .sel(IorD));
        // interfacing w/ RAM
        rw_ram IDmem 
            (.clk_100M, .clk_en, .wr_en(MemWrite), .addr(Adr), .w_data(Reg_B), .r_data(RAM_out));
        // regs for instr and data
        reg_en inst_reg
            (.clk(clk_100M), .en(IRWrite), .d(RAM_out), .q(Instr));
        reg_reset data_reg
            (.clk(clk_100M), .d(RAM_out), .q(Data));
        // instruction decoder
        ir_decode Inst_decode
            (.inst(Instr), .opcode, .funct, .rs, .rt, .rd, .shamt, .imm, .addr);
        // pre-reg file muxes
        four_mux regdest
            (.d_0(rs), .d_1(rt), .d_2(32'b11111), .d_3(32'b0), .z (Reg_A3), .sel(RegDst));
        four_mux mem_to_reg
            (.d_0(ALUOut), .d_1(Data), .d_2(PC_real), .d_3(32'b0), .z(Reg_WD3), .sel(MemtoReg));
        // interact w/ reg file
        reg_file register_file 
            (.clk(clk_100M), .wr_en(RegWrite), .w_addr(Reg_A3), .r0_addr(rs), .r1_addr(rt),
            .w_data(Reg_WD3), .r0_data(RD1_out), .r1_data(RD2_out));
        // post-register clock
        reg_reset A_reg
            (.clk(clk_100M), .d(RD1_out), .q(Reg_A));
        reg_reset B_reg
            (.clk(clk_100M), .d(RD2_out), .q(Reg_B));
        // ALUSrcA mux
        two_mux ALUSrc_A
            (.d_0(PC_real), .d_1(Reg_A), .z(SrcA), .sel(ALUSrcA));

        assign SignImm = imm[15] ? {16'b1111111111111111, imm[15:0]} : {16'b0000000000000000, imm[15:0]};
        assign Shifted_2 = SignImm << 2;
        assign shifted_addr = addr << 2;
        assign PC_first = PC_real[31:28];
        assign PCJump = {PC_first, shifted_addr};

        // ALUSrcB mux
        four_mux ALUSrc_B
            (.d_0(Reg_B), .d_1(32'b100), .d_2(SignImm), .d_3(Shifted_2), .sel(ALUSrcB), .z(SrcB));
        // run SrcA & SrcB thru ALU
        alu cpu_alu
            (.x(SrcA), .y(SrcB), .op(ALUControl), .z(ALUResult), .zero(Zero));
        // post-ALU register and mux
        reg_en result_Reg
            (.clk(clk_100M), .d(ALUResult), .q(ALUOut));
        four_mux PC_Src
            (.d_0(ALUResult), .d_1(ALUOut), .d_2(PCJump), .d_3(Reg_A), .z(PC_prime), .sel(PCSrc));

        // jump logic for BEQ and BNE
        assign PCEn = (PCWrite | (Branch & Zero) | (Branch & ~Zero));
        
endmodule
